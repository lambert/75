.TITLE SCALAR NETWORK ANALYSER - MAIN BOARD - OUTPUT STAGE - FREQUENCY RESPONSE

VS 0 1 AC 1 0 SIN(0 1 100)
C1 0 2 68p
C2 0 3 82p
C3 0 3 100p
C4 0 4 82p
C5 0 4 100p
C6 0 5 68p
C7 2 3 5.6p
C8 3 4 4.7p
C9 4 5 5.6p
L1 1 3 100nH
L2 2 4 100nH
L3 3 5 100nH
R1 0 5 50
R2 0 2 200
RS 1 2 200


.PRINT OP Iter(0) V(5)

.PRINT AC VDB(5)

*     FROM  TO  STEP
.TRAN 0     10  0.01 quiet

*       #STEPS/DECADE FROM   TO 
.AC DEC 100           100    1e9

.END
